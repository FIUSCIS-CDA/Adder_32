///////////////////////////////////////////////////////////////////////////////////
// Testbench for Component: Adder_32
// Package: FIUSCIS-CDA
// Course: CDA3102 (Computer Architecture), Florida International University
// Developer: Trevor Cickovski
// License: MIT, (C) 2020 All Rights Reserved
///////////////////////////////////////////////////////////////////////////////////


module testbench();
`include "../Test/Test.v"
///////////////////////////////////////////////////////////////////////////////////
// Inputs: A (32-bit)
//         B (32-bit)
reg[31:0] A;
reg[31:0] B;
///////////////////////////////////////////////////////////////////////////////////

///////////////////////////////////////////////////////////////////////////////////
// Outputs: S (32-bit)
wire[31:0] S;
///////////////////////////////////////////////////////////////////////////////////


Adder_32 myAdder(A, B, S);
//Test_32 myTester(S, A+B);

initial begin
////////////////////////////////////////////////////////////////////////////////////////
// Test: 45+27=72
$display("Testing: 45+27=72");
A=45; B=27;   #10;
verifyEqual32(A+B, S); 
/*if (S !== A+B) begin
           $display("Error adding %d+%d: Should be %d but got %d", A, B, A+B, S); $stop;
end*/
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: 33+142=175
$display("Testing: 33+142=175");
A=33; B=142;   #10; 
verifyEqual32(A+B, S);
/*if (S !== A+B) begin
           $display("Error adding %d+%d: Should be %d but got %d", A, B, A+B, S); $stop;
end*/
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: 0+0=0
$display("Testing: 0+0=0");
A=0; B=0;  #10;
verifyEqual32(A+B, S);
/*if (S !== A+B) begin
           $display("Error adding %d+%d: Should be %d but got %d", A, B, A+B, S); $stop;
end*/
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: -1+1=0
$display("Testing: -1+1=0");
A=-1; B=1; #10; 
verifyEqual32(A+B, S);
/*if (S !== 0) begin
           $display("Error adding %d+%d: Should be %d but got %d", A, B, 0, S); $stop;
end*/
////////////////////////////////////////////////////////////////////////////////////////

$display("All tests passed.");
end

endmodule
